module not_32(out,in);
    input [31:0] in;
    output [31:0] out;
    not not0(out[0], in[0]);
    not not1(out[1], in[1]);
    not not2(out[2], in[2]);
    not not3(out[3], in[3]);
    not not4(out[4], in[4]);
    not not5(out[5], in[5]);
    not not6(out[6], in[6]);
    not not7(out[7], in[7]);
    not not8(out[8], in[8]);
    not not9(out[9], in[9]);
    not not10(out[10], in[10]);
    not not11(out[11], in[11]);
    not not12(out[12], in[12]);
    not not13(out[13], in[13]);
    not not14(out[14], in[14]);
    not not15(out[15], in[15]);
    not not16(out[16], in[16]);
    not not17(out[17], in[17]);
    not not18(out[18], in[18]);
    not not19(out[19], in[19]);
    not not20(out[20], in[20]);
    not not21(out[21], in[21]);
    not not22(out[22], in[22]);
    not not23(out[23], in[23]);
    not not24(out[24], in[24]);
    not not25(out[25], in[25]);
    not not26(out[26], in[26]);
    not not27(out[27], in[27]);
    not not28(out[28], in[28]);
    not not29(out[29], in[29]);
    not not30(out[30], in[30]);
    not not31(out[31], in[31]);
endmodule